-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity SDRAMTest_ROM is
generic
	(
		maxAddrBit : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end SDRAMTest_ROM;

architecture arch of SDRAMTest_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBit+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0ba08080",
     1 => x"df040000",
     2 => x"80047004",
     3 => x"71fd0608",
     4 => x"72830609",
     5 => x"81058205",
     6 => x"832b2a83",
     7 => x"ffff0652",
     8 => x"0471fc06",
     9 => x"08728306",
    10 => x"09810583",
    11 => x"05101010",
    12 => x"2a81ff06",
    13 => x"520471fc",
    14 => x"06080ba0",
    15 => x"808cc873",
    16 => x"83061010",
    17 => x"05080673",
    18 => x"81ff0673",
    19 => x"83060981",
    20 => x"05830510",
    21 => x"10102b07",
    22 => x"72fc060c",
    23 => x"5151040b",
    24 => x"a08080ea",
    25 => x"0ba0808b",
    26 => x"c5040ba0",
    27 => x"8080ea04",
    28 => x"00000002",
    29 => x"f8050d73",
    30 => x"52ff8408",
    31 => x"70882a70",
    32 => x"81065151",
    33 => x"5170802e",
    34 => x"f03871ff",
    35 => x"840c71a0",
    36 => x"8092d80c",
    37 => x"0288050d",
    38 => x"0402f005",
    39 => x"0d755380",
    40 => x"73337081",
    41 => x"ff065353",
    42 => x"5470742e",
    43 => x"ac387181",
    44 => x"ff068114",
    45 => x"5452ff84",
    46 => x"0870882a",
    47 => x"70810651",
    48 => x"51517080",
    49 => x"2ef03871",
    50 => x"ff840c81",
    51 => x"14733370",
    52 => x"81ff0653",
    53 => x"535470d6",
    54 => x"3873a080",
    55 => x"92d80c02",
    56 => x"90050d04",
    57 => x"02c4050d",
    58 => x"0280c005",
    59 => x"a08093b8",
    60 => x"5b568076",
    61 => x"70840558",
    62 => x"08715e5e",
    63 => x"577c7084",
    64 => x"055e0858",
    65 => x"805b7798",
    66 => x"2a78882b",
    67 => x"59537288",
    68 => x"38765ea0",
    69 => x"80848904",
    70 => x"7b802e81",
    71 => x"c638805c",
    72 => x"7280e42e",
    73 => x"9f387280",
    74 => x"e4268d38",
    75 => x"7280e32e",
    76 => x"80ee38a0",
    77 => x"8083ad04",
    78 => x"7280f32e",
    79 => x"80cc38a0",
    80 => x"8083ad04",
    81 => x"75841771",
    82 => x"087e5c56",
    83 => x"57528755",
    84 => x"739c2a74",
    85 => x"842b5552",
    86 => x"71802e83",
    87 => x"38815989",
    88 => x"72258938",
    89 => x"b71252a0",
    90 => x"8082ef04",
    91 => x"b0125278",
    92 => x"802e8838",
    93 => x"7151a080",
    94 => x"80f32dff",
    95 => x"15557480",
    96 => x"25ce3880",
    97 => x"54a08083",
    98 => x"c3047584",
    99 => x"17710870",
   100 => x"545c5752",
   101 => x"a0808199",
   102 => x"2d7b54a0",
   103 => x"8083c304",
   104 => x"75841771",
   105 => x"08555752",
   106 => x"a08083f2",
   107 => x"04a551a0",
   108 => x"8080f32d",
   109 => x"7251a080",
   110 => x"80f32d82",
   111 => x"1757a080",
   112 => x"83fc0473",
   113 => x"ff155552",
   114 => x"807225b0",
   115 => x"38797081",
   116 => x"055b3370",
   117 => x"5253a080",
   118 => x"80f32d81",
   119 => x"1757a080",
   120 => x"83c30472",
   121 => x"a52e0981",
   122 => x"06883881",
   123 => x"5ca08083",
   124 => x"fc047251",
   125 => x"a08080f3",
   126 => x"2d811757",
   127 => x"811b5b83",
   128 => x"7b25fe82",
   129 => x"3872fdf5",
   130 => x"387da080",
   131 => x"92d80c02",
   132 => x"bc050d04",
   133 => x"02f4050d",
   134 => x"74765253",
   135 => x"80712590",
   136 => x"38705272",
   137 => x"70840554",
   138 => x"08ff1353",
   139 => x"5171f438",
   140 => x"028c050d",
   141 => x"0402d805",
   142 => x"0d7b7d5b",
   143 => x"56810ba0",
   144 => x"808cd859",
   145 => x"57835977",
   146 => x"08760c75",
   147 => x"08780856",
   148 => x"5473752e",
   149 => x"92387508",
   150 => x"537452a0",
   151 => x"808ce851",
   152 => x"a08081e4",
   153 => x"2d805779",
   154 => x"527551a0",
   155 => x"8084942d",
   156 => x"75085473",
   157 => x"752e9238",
   158 => x"75085374",
   159 => x"52a0808d",
   160 => x"a851a080",
   161 => x"81e42d80",
   162 => x"57ff1984",
   163 => x"19595978",
   164 => x"8025ffb3",
   165 => x"3876a080",
   166 => x"92d80c02",
   167 => x"a8050d04",
   168 => x"02ec050d",
   169 => x"76548155",
   170 => x"85aad5aa",
   171 => x"d5740cfa",
   172 => x"d5aad5aa",
   173 => x"0b8c150c",
   174 => x"cc7434b3",
   175 => x"0b8f1534",
   176 => x"73085372",
   177 => x"fce2d5aa",
   178 => x"d52e9038",
   179 => x"730852a0",
   180 => x"808de851",
   181 => x"a08081e4",
   182 => x"2d80558c",
   183 => x"14085372",
   184 => x"fad5aad4",
   185 => x"b32e9138",
   186 => x"8c140852",
   187 => x"a0808ea4",
   188 => x"51a08081",
   189 => x"e42d8055",
   190 => x"77527351",
   191 => x"a0808494",
   192 => x"2d730853",
   193 => x"72fce2d5",
   194 => x"aad52e90",
   195 => x"38730852",
   196 => x"a0808ee0",
   197 => x"51a08081",
   198 => x"e42d8055",
   199 => x"8c140853",
   200 => x"72fad5aa",
   201 => x"d4b32e91",
   202 => x"388c1408",
   203 => x"52a0808f",
   204 => x"9c51a080",
   205 => x"81e42d80",
   206 => x"5574a080",
   207 => x"92d80c02",
   208 => x"94050d04",
   209 => x"02c8050d",
   210 => x"7f5c800b",
   211 => x"a0808fd8",
   212 => x"525ba080",
   213 => x"81e42d80",
   214 => x"e1b3578e",
   215 => x"5d76598f",
   216 => x"ffff5a76",
   217 => x"bfffff06",
   218 => x"77107096",
   219 => x"2a708106",
   220 => x"51575858",
   221 => x"74802e85",
   222 => x"38768107",
   223 => x"5776952a",
   224 => x"70810651",
   225 => x"5574802e",
   226 => x"85387681",
   227 => x"325776bf",
   228 => x"ffff0678",
   229 => x"84291d79",
   230 => x"710c5670",
   231 => x"84291d56",
   232 => x"750c7610",
   233 => x"70962a70",
   234 => x"81065156",
   235 => x"5774802e",
   236 => x"85387681",
   237 => x"07577695",
   238 => x"2a708106",
   239 => x"51557480",
   240 => x"2e853876",
   241 => x"813257ff",
   242 => x"1a5a7980",
   243 => x"25ff9438",
   244 => x"78578fff",
   245 => x"ff5a76bf",
   246 => x"ffff0677",
   247 => x"1070962a",
   248 => x"70810651",
   249 => x"57585674",
   250 => x"802e8538",
   251 => x"76810757",
   252 => x"76952a70",
   253 => x"81065155",
   254 => x"74802e85",
   255 => x"38768132",
   256 => x"5776bfff",
   257 => x"ff067684",
   258 => x"291d7008",
   259 => x"7284291f",
   260 => x"70085152",
   261 => x"5b565878",
   262 => x"762ea638",
   263 => x"807b53a0",
   264 => x"808fec52",
   265 => x"5ea08081",
   266 => x"e42d7854",
   267 => x"75537552",
   268 => x"a0809080",
   269 => x"51a08081",
   270 => x"e42d7d5b",
   271 => x"a08088c4",
   272 => x"04811b5b",
   273 => x"74782ea6",
   274 => x"38807b53",
   275 => x"a0808fec",
   276 => x"525ea080",
   277 => x"81e42d74",
   278 => x"54775377",
   279 => x"52a08090",
   280 => x"8051a080",
   281 => x"81e42d7d",
   282 => x"5ba08088",
   283 => x"f104811b",
   284 => x"5b761070",
   285 => x"962a7081",
   286 => x"06515657",
   287 => x"74802e85",
   288 => x"38768107",
   289 => x"5776952a",
   290 => x"70810651",
   291 => x"5574802e",
   292 => x"85387681",
   293 => x"3257ff1a",
   294 => x"5a798025",
   295 => x"feb838ff",
   296 => x"1d5d7cfd",
   297 => x"b8387da0",
   298 => x"8092d80c",
   299 => x"02b8050d",
   300 => x"0402d005",
   301 => x"0d7d5b81",
   302 => x"5a805980",
   303 => x"c07a595c",
   304 => x"85ada989",
   305 => x"bb7b0c79",
   306 => x"57815697",
   307 => x"55777607",
   308 => x"822b7b11",
   309 => x"515485ad",
   310 => x"a989bb74",
   311 => x"0c7510ff",
   312 => x"16565674",
   313 => x"8025e638",
   314 => x"77108118",
   315 => x"58589877",
   316 => x"25d7387e",
   317 => x"527a51a0",
   318 => x"8084942d",
   319 => x"8158ff87",
   320 => x"87a5c37b",
   321 => x"0c975777",
   322 => x"822b7b11",
   323 => x"70085656",
   324 => x"5673ff87",
   325 => x"87a5c32e",
   326 => x"0981068a",
   327 => x"38787807",
   328 => x"59a0808a",
   329 => x"c3047408",
   330 => x"547385ad",
   331 => x"a989bb2e",
   332 => x"92388075",
   333 => x"08547653",
   334 => x"a08090a8",
   335 => x"525aa080",
   336 => x"81e42d77",
   337 => x"10ff1858",
   338 => x"58768025",
   339 => x"ffb93878",
   340 => x"822b5978",
   341 => x"802eb838",
   342 => x"7852a080",
   343 => x"90c851a0",
   344 => x"8081e42d",
   345 => x"78992a81",
   346 => x"32708106",
   347 => x"70098105",
   348 => x"70720770",
   349 => x"09709f2c",
   350 => x"7f067e10",
   351 => x"87fffffe",
   352 => x"0662812c",
   353 => x"435f5f51",
   354 => x"51565155",
   355 => x"78d63879",
   356 => x"09810570",
   357 => x"7b079f2a",
   358 => x"51547bbf",
   359 => x"24903873",
   360 => x"802e8b38",
   361 => x"a08090e0",
   362 => x"51a08081",
   363 => x"e42d7b52",
   364 => x"a08091ac",
   365 => x"51a08081",
   366 => x"e42d79a0",
   367 => x"8092d80c",
   368 => x"02b0050d",
   369 => x"0402f805",
   370 => x"0d88bd0b",
   371 => x"ff880ca0",
   372 => x"80528051",
   373 => x"a08084b5",
   374 => x"2da08092",
   375 => x"d808802e",
   376 => x"8b38a080",
   377 => x"91e851a0",
   378 => x"8081e42d",
   379 => x"a0805280",
   380 => x"51a08085",
   381 => x"a02da080",
   382 => x"92d80880",
   383 => x"2e8b38a0",
   384 => x"80928c51",
   385 => x"a08081e4",
   386 => x"2da08052",
   387 => x"8051a080",
   388 => x"89b12da0",
   389 => x"8092d808",
   390 => x"802e8b38",
   391 => x"a08092a8",
   392 => x"51a08081",
   393 => x"e42d8051",
   394 => x"a08086c4",
   395 => x"2da08092",
   396 => x"d808802e",
   397 => x"ff9938a0",
   398 => x"8092c051",
   399 => x"a08081e4",
   400 => x"2da0808b",
   401 => x"cf040000",
   402 => x"00ffffff",
   403 => x"ff00ffff",
   404 => x"ffff00ff",
   405 => x"ffffff00",
   406 => x"00000000",
   407 => x"55555555",
   408 => x"aaaaaaaa",
   409 => x"ffffffff",
   410 => x"53616e69",
   411 => x"74792063",
   412 => x"6865636b",
   413 => x"20666169",
   414 => x"6c656420",
   415 => x"28626566",
   416 => x"6f726520",
   417 => x"63616368",
   418 => x"65207265",
   419 => x"66726573",
   420 => x"6829206f",
   421 => x"6e203078",
   422 => x"25642028",
   423 => x"676f7420",
   424 => x"30782564",
   425 => x"290a0000",
   426 => x"53616e69",
   427 => x"74792063",
   428 => x"6865636b",
   429 => x"20666169",
   430 => x"6c656420",
   431 => x"28616674",
   432 => x"65722063",
   433 => x"61636865",
   434 => x"20726566",
   435 => x"72657368",
   436 => x"29206f6e",
   437 => x"20307825",
   438 => x"64202867",
   439 => x"6f742030",
   440 => x"78256429",
   441 => x"0a000000",
   442 => x"42797465",
   443 => x"20636865",
   444 => x"636b2066",
   445 => x"61696c65",
   446 => x"64202862",
   447 => x"65666f72",
   448 => x"65206361",
   449 => x"63686520",
   450 => x"72656672",
   451 => x"65736829",
   452 => x"20617420",
   453 => x"30202867",
   454 => x"6f742030",
   455 => x"78256429",
   456 => x"0a000000",
   457 => x"42797465",
   458 => x"20636865",
   459 => x"636b2066",
   460 => x"61696c65",
   461 => x"64202862",
   462 => x"65666f72",
   463 => x"65206361",
   464 => x"63686520",
   465 => x"72656672",
   466 => x"65736829",
   467 => x"20617420",
   468 => x"33202867",
   469 => x"6f742030",
   470 => x"78256429",
   471 => x"0a000000",
   472 => x"42797465",
   473 => x"20636865",
   474 => x"636b2066",
   475 => x"61696c65",
   476 => x"64202861",
   477 => x"66746572",
   478 => x"20636163",
   479 => x"68652072",
   480 => x"65667265",
   481 => x"73682920",
   482 => x"61742030",
   483 => x"2028676f",
   484 => x"74203078",
   485 => x"2564290a",
   486 => x"00000000",
   487 => x"42797465",
   488 => x"20636865",
   489 => x"636b2066",
   490 => x"61696c65",
   491 => x"64202861",
   492 => x"66746572",
   493 => x"20636163",
   494 => x"68652072",
   495 => x"65667265",
   496 => x"73682920",
   497 => x"61742033",
   498 => x"2028676f",
   499 => x"74203078",
   500 => x"2564290a",
   501 => x"00000000",
   502 => x"43686563",
   503 => x"6b696e67",
   504 => x"206d656d",
   505 => x"6f72792e",
   506 => x"2e2e0a00",
   507 => x"30782564",
   508 => x"20676f6f",
   509 => x"64207265",
   510 => x"6164732c",
   511 => x"20000000",
   512 => x"4572726f",
   513 => x"72206174",
   514 => x"20307825",
   515 => x"642c2065",
   516 => x"78706563",
   517 => x"74656420",
   518 => x"30782564",
   519 => x"2c20676f",
   520 => x"74203078",
   521 => x"25640a00",
   522 => x"42616420",
   523 => x"64617461",
   524 => x"20666f75",
   525 => x"6e642061",
   526 => x"74203078",
   527 => x"25642028",
   528 => x"30782564",
   529 => x"290a0000",
   530 => x"416c6961",
   531 => x"73657320",
   532 => x"666f756e",
   533 => x"64206174",
   534 => x"20307825",
   535 => x"640a0000",
   536 => x"28416c69",
   537 => x"61736573",
   538 => x"2070726f",
   539 => x"6261626c",
   540 => x"79207369",
   541 => x"6d706c79",
   542 => x"20696e64",
   543 => x"69636174",
   544 => x"65207468",
   545 => x"61742052",
   546 => x"414d0a69",
   547 => x"7320736d",
   548 => x"616c6c65",
   549 => x"72207468",
   550 => x"616e2036",
   551 => x"34206d65",
   552 => x"67616279",
   553 => x"74657329",
   554 => x"0a000000",
   555 => x"53445241",
   556 => x"4d207369",
   557 => x"7a652028",
   558 => x"61737375",
   559 => x"6d696e67",
   560 => x"206e6f20",
   561 => x"61646472",
   562 => x"65737320",
   563 => x"6661756c",
   564 => x"74732920",
   565 => x"69732030",
   566 => x"78256420",
   567 => x"6d656761",
   568 => x"62797465",
   569 => x"730a0000",
   570 => x"46697273",
   571 => x"74207374",
   572 => x"61676520",
   573 => x"73616e69",
   574 => x"74792063",
   575 => x"6865636b",
   576 => x"20706173",
   577 => x"7365642e",
   578 => x"0a000000",
   579 => x"42797465",
   580 => x"20286471",
   581 => x"6d292063",
   582 => x"6865636b",
   583 => x"20706173",
   584 => x"7365640a",
   585 => x"00000000",
   586 => x"41646472",
   587 => x"65737320",
   588 => x"63686563",
   589 => x"6b207061",
   590 => x"73736564",
   591 => x"2e0a0000",
   592 => x"4c465352",
   593 => x"20636865",
   594 => x"636b2070",
   595 => x"61737365",
   596 => x"642e0a0a",
   597 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBit-1 downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBit-1 downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr)));
		end if;
	end if;
end process;


end arch;

