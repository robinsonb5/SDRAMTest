-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity SDRAMTest_ROM is
generic
	(
		maxAddrBit : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end SDRAMTest_ROM;

architecture arch of SDRAMTest_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBit+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0ba08080",
     1 => x"df040000",
     2 => x"80047004",
     3 => x"71fd0608",
     4 => x"72830609",
     5 => x"81058205",
     6 => x"832b2a83",
     7 => x"ffff0652",
     8 => x"0471fc06",
     9 => x"08728306",
    10 => x"09810583",
    11 => x"05101010",
    12 => x"2a81ff06",
    13 => x"520471fc",
    14 => x"06080ba0",
    15 => x"808cdc73",
    16 => x"83061010",
    17 => x"05080673",
    18 => x"81ff0673",
    19 => x"83060981",
    20 => x"05830510",
    21 => x"10102b07",
    22 => x"72fc060c",
    23 => x"5151040b",
    24 => x"a08080ea",
    25 => x"0ba0808b",
    26 => x"d9040ba0",
    27 => x"8080ea04",
    28 => x"00000002",
    29 => x"f8050d73",
    30 => x"52ff8408",
    31 => x"70882a70",
    32 => x"81065151",
    33 => x"5170802e",
    34 => x"f03871ff",
    35 => x"840c71a0",
    36 => x"8092ec0c",
    37 => x"0288050d",
    38 => x"0402f005",
    39 => x"0d755380",
    40 => x"73a08080",
    41 => x"a12d7081",
    42 => x"ff065353",
    43 => x"5470742e",
    44 => x"b0387181",
    45 => x"ff068114",
    46 => x"5452ff84",
    47 => x"0870882a",
    48 => x"70810651",
    49 => x"51517080",
    50 => x"2ef03871",
    51 => x"ff840c81",
    52 => x"1473a080",
    53 => x"80a12d70",
    54 => x"81ff0653",
    55 => x"535470d2",
    56 => x"3873a080",
    57 => x"92ec0c02",
    58 => x"90050d04",
    59 => x"02c4050d",
    60 => x"0280c005",
    61 => x"a08093cc",
    62 => x"5b568076",
    63 => x"70840558",
    64 => x"08715e5e",
    65 => x"577c7084",
    66 => x"055e0858",
    67 => x"805b7798",
    68 => x"2a78882b",
    69 => x"59537288",
    70 => x"38765ea0",
    71 => x"80849504",
    72 => x"7b802e81",
    73 => x"ca38805c",
    74 => x"7280e42e",
    75 => x"9f387280",
    76 => x"e4268d38",
    77 => x"7280e32e",
    78 => x"80ee38a0",
    79 => x"8083b504",
    80 => x"7280f32e",
    81 => x"80cc38a0",
    82 => x"8083b504",
    83 => x"75841771",
    84 => x"087e5c56",
    85 => x"57528755",
    86 => x"739c2a74",
    87 => x"842b5552",
    88 => x"71802e83",
    89 => x"38815989",
    90 => x"72258938",
    91 => x"b71252a0",
    92 => x"8082f704",
    93 => x"b0125278",
    94 => x"802e8838",
    95 => x"7151a080",
    96 => x"80f32dff",
    97 => x"15557480",
    98 => x"25ce3880",
    99 => x"54a08083",
   100 => x"cb047584",
   101 => x"17710870",
   102 => x"545c5752",
   103 => x"a0808199",
   104 => x"2d7b54a0",
   105 => x"8083cb04",
   106 => x"75841771",
   107 => x"08555752",
   108 => x"a08083fe",
   109 => x"04a551a0",
   110 => x"8080f32d",
   111 => x"7251a080",
   112 => x"80f32d82",
   113 => x"1757a080",
   114 => x"84880473",
   115 => x"ff155552",
   116 => x"807225b4",
   117 => x"38797081",
   118 => x"055ba080",
   119 => x"80a12d70",
   120 => x"5253a080",
   121 => x"80f32d81",
   122 => x"1757a080",
   123 => x"83cb0472",
   124 => x"a52e0981",
   125 => x"06883881",
   126 => x"5ca08084",
   127 => x"88047251",
   128 => x"a08080f3",
   129 => x"2d811757",
   130 => x"811b5b83",
   131 => x"7b25fdfe",
   132 => x"3872fdf1",
   133 => x"387da080",
   134 => x"92ec0c02",
   135 => x"bc050d04",
   136 => x"02f4050d",
   137 => x"74765253",
   138 => x"80712590",
   139 => x"38705272",
   140 => x"70840554",
   141 => x"08ff1353",
   142 => x"5171f438",
   143 => x"028c050d",
   144 => x"0402d805",
   145 => x"0d7b7d5b",
   146 => x"56810ba0",
   147 => x"808cec59",
   148 => x"57835977",
   149 => x"08760c75",
   150 => x"08780856",
   151 => x"5473752e",
   152 => x"92387508",
   153 => x"537452a0",
   154 => x"808cfc51",
   155 => x"a08081ec",
   156 => x"2d805779",
   157 => x"527551a0",
   158 => x"8084a02d",
   159 => x"75085473",
   160 => x"752e9238",
   161 => x"75085374",
   162 => x"52a0808d",
   163 => x"bc51a080",
   164 => x"81ec2d80",
   165 => x"57ff1984",
   166 => x"19595978",
   167 => x"8025ffb3",
   168 => x"3876a080",
   169 => x"92ec0c02",
   170 => x"a8050d04",
   171 => x"02ec050d",
   172 => x"76548155",
   173 => x"85aad5aa",
   174 => x"d5740cfa",
   175 => x"d5aad5aa",
   176 => x"0b8c150c",
   177 => x"cc74a080",
   178 => x"80b62db3",
   179 => x"0b8f15a0",
   180 => x"8080b62d",
   181 => x"73085372",
   182 => x"fce2d5aa",
   183 => x"d52e9038",
   184 => x"730852a0",
   185 => x"808dfc51",
   186 => x"a08081ec",
   187 => x"2d80558c",
   188 => x"14085372",
   189 => x"fad5aad4",
   190 => x"b32e9138",
   191 => x"8c140852",
   192 => x"a0808eb8",
   193 => x"51a08081",
   194 => x"ec2d8055",
   195 => x"77527351",
   196 => x"a08084a0",
   197 => x"2d730853",
   198 => x"72fce2d5",
   199 => x"aad52e90",
   200 => x"38730852",
   201 => x"a0808ef4",
   202 => x"51a08081",
   203 => x"ec2d8055",
   204 => x"8c140853",
   205 => x"72fad5aa",
   206 => x"d4b32e91",
   207 => x"388c1408",
   208 => x"52a0808f",
   209 => x"b051a080",
   210 => x"81ec2d80",
   211 => x"5574a080",
   212 => x"92ec0c02",
   213 => x"94050d04",
   214 => x"02c8050d",
   215 => x"7f5c800b",
   216 => x"a0808fec",
   217 => x"525ba080",
   218 => x"81ec2d80",
   219 => x"e1b3578e",
   220 => x"5d76598f",
   221 => x"ffff5a76",
   222 => x"bfffff06",
   223 => x"77107096",
   224 => x"2a708106",
   225 => x"51575858",
   226 => x"74802e85",
   227 => x"38768107",
   228 => x"5776952a",
   229 => x"70810651",
   230 => x"5574802e",
   231 => x"85387681",
   232 => x"325776bf",
   233 => x"ffff0678",
   234 => x"84291d79",
   235 => x"710c5670",
   236 => x"84291d56",
   237 => x"750c7610",
   238 => x"70962a70",
   239 => x"81065156",
   240 => x"5774802e",
   241 => x"85387681",
   242 => x"07577695",
   243 => x"2a708106",
   244 => x"51557480",
   245 => x"2e853876",
   246 => x"813257ff",
   247 => x"1a5a7980",
   248 => x"25ff9438",
   249 => x"78578fff",
   250 => x"ff5a76bf",
   251 => x"ffff0677",
   252 => x"1070962a",
   253 => x"70810651",
   254 => x"57585674",
   255 => x"802e8538",
   256 => x"76810757",
   257 => x"76952a70",
   258 => x"81065155",
   259 => x"74802e85",
   260 => x"38768132",
   261 => x"5776bfff",
   262 => x"ff067684",
   263 => x"291d7008",
   264 => x"7284291f",
   265 => x"70085152",
   266 => x"5b565878",
   267 => x"762ea638",
   268 => x"807b53a0",
   269 => x"80908052",
   270 => x"5ea08081",
   271 => x"ec2d7854",
   272 => x"75537552",
   273 => x"a0809094",
   274 => x"51a08081",
   275 => x"ec2d7d5b",
   276 => x"a08088d8",
   277 => x"04811b5b",
   278 => x"74782ea6",
   279 => x"38807b53",
   280 => x"a0809080",
   281 => x"525ea080",
   282 => x"81ec2d74",
   283 => x"54775377",
   284 => x"52a08090",
   285 => x"9451a080",
   286 => x"81ec2d7d",
   287 => x"5ba08089",
   288 => x"8504811b",
   289 => x"5b761070",
   290 => x"962a7081",
   291 => x"06515657",
   292 => x"74802e85",
   293 => x"38768107",
   294 => x"5776952a",
   295 => x"70810651",
   296 => x"5574802e",
   297 => x"85387681",
   298 => x"3257ff1a",
   299 => x"5a798025",
   300 => x"feb838ff",
   301 => x"1d5d7cfd",
   302 => x"b8387da0",
   303 => x"8092ec0c",
   304 => x"02b8050d",
   305 => x"0402d005",
   306 => x"0d7d5b81",
   307 => x"5a805980",
   308 => x"c07a595c",
   309 => x"85ada989",
   310 => x"bb7b0c79",
   311 => x"57815697",
   312 => x"55777607",
   313 => x"822b7b11",
   314 => x"515485ad",
   315 => x"a989bb74",
   316 => x"0c7510ff",
   317 => x"16565674",
   318 => x"8025e638",
   319 => x"77108118",
   320 => x"58589877",
   321 => x"25d7387e",
   322 => x"527a51a0",
   323 => x"8084a02d",
   324 => x"8158ff87",
   325 => x"87a5c37b",
   326 => x"0c975777",
   327 => x"822b7b11",
   328 => x"70085656",
   329 => x"5673ff87",
   330 => x"87a5c32e",
   331 => x"0981068a",
   332 => x"38787807",
   333 => x"59a0808a",
   334 => x"d7047408",
   335 => x"547385ad",
   336 => x"a989bb2e",
   337 => x"92388075",
   338 => x"08547653",
   339 => x"a08090bc",
   340 => x"525aa080",
   341 => x"81ec2d77",
   342 => x"10ff1858",
   343 => x"58768025",
   344 => x"ffb93878",
   345 => x"822b5978",
   346 => x"802eb838",
   347 => x"7852a080",
   348 => x"90dc51a0",
   349 => x"8081ec2d",
   350 => x"78992a81",
   351 => x"32708106",
   352 => x"70098105",
   353 => x"70720770",
   354 => x"09709f2c",
   355 => x"7f067e10",
   356 => x"87fffffe",
   357 => x"0662812c",
   358 => x"435f5f51",
   359 => x"51565155",
   360 => x"78d63879",
   361 => x"09810570",
   362 => x"7b079f2a",
   363 => x"51547bbf",
   364 => x"24903873",
   365 => x"802e8b38",
   366 => x"a08090f4",
   367 => x"51a08081",
   368 => x"ec2d7b52",
   369 => x"a08091c0",
   370 => x"51a08081",
   371 => x"ec2d79a0",
   372 => x"8092ec0c",
   373 => x"02b0050d",
   374 => x"0402f805",
   375 => x"0d88bd0b",
   376 => x"ff880ca0",
   377 => x"80528051",
   378 => x"a08084c1",
   379 => x"2da08092",
   380 => x"ec08802e",
   381 => x"8b38a080",
   382 => x"91fc51a0",
   383 => x"8081ec2d",
   384 => x"a0805280",
   385 => x"51a08085",
   386 => x"ac2da080",
   387 => x"92ec0880",
   388 => x"2e8b38a0",
   389 => x"8092a051",
   390 => x"a08081ec",
   391 => x"2da08052",
   392 => x"8051a080",
   393 => x"89c52da0",
   394 => x"8092ec08",
   395 => x"802e8b38",
   396 => x"a08092bc",
   397 => x"51a08081",
   398 => x"ec2d8051",
   399 => x"a08086d8",
   400 => x"2da08092",
   401 => x"ec08802e",
   402 => x"ff9938a0",
   403 => x"8092d451",
   404 => x"a08081ec",
   405 => x"2da0808b",
   406 => x"e3040000",
   407 => x"00ffffff",
   408 => x"ff00ffff",
   409 => x"ffff00ff",
   410 => x"ffffff00",
   411 => x"00000000",
   412 => x"55555555",
   413 => x"aaaaaaaa",
   414 => x"ffffffff",
   415 => x"53616e69",
   416 => x"74792063",
   417 => x"6865636b",
   418 => x"20666169",
   419 => x"6c656420",
   420 => x"28626566",
   421 => x"6f726520",
   422 => x"63616368",
   423 => x"65207265",
   424 => x"66726573",
   425 => x"6829206f",
   426 => x"6e203078",
   427 => x"25642028",
   428 => x"676f7420",
   429 => x"30782564",
   430 => x"290a0000",
   431 => x"53616e69",
   432 => x"74792063",
   433 => x"6865636b",
   434 => x"20666169",
   435 => x"6c656420",
   436 => x"28616674",
   437 => x"65722063",
   438 => x"61636865",
   439 => x"20726566",
   440 => x"72657368",
   441 => x"29206f6e",
   442 => x"20307825",
   443 => x"64202867",
   444 => x"6f742030",
   445 => x"78256429",
   446 => x"0a000000",
   447 => x"42797465",
   448 => x"20636865",
   449 => x"636b2066",
   450 => x"61696c65",
   451 => x"64202862",
   452 => x"65666f72",
   453 => x"65206361",
   454 => x"63686520",
   455 => x"72656672",
   456 => x"65736829",
   457 => x"20617420",
   458 => x"30202867",
   459 => x"6f742030",
   460 => x"78256429",
   461 => x"0a000000",
   462 => x"42797465",
   463 => x"20636865",
   464 => x"636b2066",
   465 => x"61696c65",
   466 => x"64202862",
   467 => x"65666f72",
   468 => x"65206361",
   469 => x"63686520",
   470 => x"72656672",
   471 => x"65736829",
   472 => x"20617420",
   473 => x"33202867",
   474 => x"6f742030",
   475 => x"78256429",
   476 => x"0a000000",
   477 => x"42797465",
   478 => x"20636865",
   479 => x"636b2066",
   480 => x"61696c65",
   481 => x"64202861",
   482 => x"66746572",
   483 => x"20636163",
   484 => x"68652072",
   485 => x"65667265",
   486 => x"73682920",
   487 => x"61742030",
   488 => x"2028676f",
   489 => x"74203078",
   490 => x"2564290a",
   491 => x"00000000",
   492 => x"42797465",
   493 => x"20636865",
   494 => x"636b2066",
   495 => x"61696c65",
   496 => x"64202861",
   497 => x"66746572",
   498 => x"20636163",
   499 => x"68652072",
   500 => x"65667265",
   501 => x"73682920",
   502 => x"61742033",
   503 => x"2028676f",
   504 => x"74203078",
   505 => x"2564290a",
   506 => x"00000000",
   507 => x"43686563",
   508 => x"6b696e67",
   509 => x"206d656d",
   510 => x"6f72792e",
   511 => x"2e2e0a00",
   512 => x"30782564",
   513 => x"20676f6f",
   514 => x"64207265",
   515 => x"6164732c",
   516 => x"20000000",
   517 => x"4572726f",
   518 => x"72206174",
   519 => x"20307825",
   520 => x"642c2065",
   521 => x"78706563",
   522 => x"74656420",
   523 => x"30782564",
   524 => x"2c20676f",
   525 => x"74203078",
   526 => x"25640a00",
   527 => x"42616420",
   528 => x"64617461",
   529 => x"20666f75",
   530 => x"6e642061",
   531 => x"74203078",
   532 => x"25642028",
   533 => x"30782564",
   534 => x"290a0000",
   535 => x"416c6961",
   536 => x"73657320",
   537 => x"666f756e",
   538 => x"64206174",
   539 => x"20307825",
   540 => x"640a0000",
   541 => x"28416c69",
   542 => x"61736573",
   543 => x"2070726f",
   544 => x"6261626c",
   545 => x"79207369",
   546 => x"6d706c79",
   547 => x"20696e64",
   548 => x"69636174",
   549 => x"65207468",
   550 => x"61742052",
   551 => x"414d0a69",
   552 => x"7320736d",
   553 => x"616c6c65",
   554 => x"72207468",
   555 => x"616e2036",
   556 => x"34206d65",
   557 => x"67616279",
   558 => x"74657329",
   559 => x"0a000000",
   560 => x"53445241",
   561 => x"4d207369",
   562 => x"7a652028",
   563 => x"61737375",
   564 => x"6d696e67",
   565 => x"206e6f20",
   566 => x"61646472",
   567 => x"65737320",
   568 => x"6661756c",
   569 => x"74732920",
   570 => x"69732030",
   571 => x"78256420",
   572 => x"6d656761",
   573 => x"62797465",
   574 => x"730a0000",
   575 => x"46697273",
   576 => x"74207374",
   577 => x"61676520",
   578 => x"73616e69",
   579 => x"74792063",
   580 => x"6865636b",
   581 => x"20706173",
   582 => x"7365642e",
   583 => x"0a000000",
   584 => x"42797465",
   585 => x"20286471",
   586 => x"6d292063",
   587 => x"6865636b",
   588 => x"20706173",
   589 => x"7365640a",
   590 => x"00000000",
   591 => x"41646472",
   592 => x"65737320",
   593 => x"63686563",
   594 => x"6b207061",
   595 => x"73736564",
   596 => x"2e0a0000",
   597 => x"4c465352",
   598 => x"20636865",
   599 => x"636b2070",
   600 => x"61737365",
   601 => x"642e0a0a",
   602 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBit downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBit downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBit downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBit downto 2))));
		end if;
	end if;
end process;


end arch;

