-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity SDRAMTest_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end SDRAMTest_ROM;

architecture arch of SDRAMTest_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"84808080",
     1 => x"ed040000",
     2 => x"00000000",
     3 => x"84808080",
     4 => x"880d8004",
     5 => x"84808080",
     6 => x"940471fd",
     7 => x"06087283",
     8 => x"06098105",
     9 => x"8205832b",
    10 => x"2a83ffff",
    11 => x"06520471",
    12 => x"fc060872",
    13 => x"83060981",
    14 => x"05830510",
    15 => x"10102a81",
    16 => x"ff065204",
    17 => x"71fc0608",
    18 => x"8480808d",
    19 => x"84738306",
    20 => x"10100508",
    21 => x"067381ff",
    22 => x"06738306",
    23 => x"09810583",
    24 => x"05101010",
    25 => x"2b0772fc",
    26 => x"060c5151",
    27 => x"04028405",
    28 => x"84808080",
    29 => x"880c8480",
    30 => x"8080940b",
    31 => x"8480808b",
    32 => x"e7040000",
    33 => x"02f8050d",
    34 => x"7352ff84",
    35 => x"0870882a",
    36 => x"70810651",
    37 => x"51517080",
    38 => x"2ef03871",
    39 => x"ff840c71",
    40 => x"84808093",
    41 => x"900c0288",
    42 => x"050d0402",
    43 => x"f0050d75",
    44 => x"53807384",
    45 => x"808080af",
    46 => x"2d7081ff",
    47 => x"06535354",
    48 => x"70742eb1",
    49 => x"387181ff",
    50 => x"06811454",
    51 => x"52ff8408",
    52 => x"70882a70",
    53 => x"81065151",
    54 => x"5170802e",
    55 => x"f03871ff",
    56 => x"840c8114",
    57 => x"73848080",
    58 => x"80af2d70",
    59 => x"81ff0653",
    60 => x"535470d1",
    61 => x"38738480",
    62 => x"8093900c",
    63 => x"0290050d",
    64 => x"0402c405",
    65 => x"0d0280c0",
    66 => x"05848080",
    67 => x"93f05b56",
    68 => x"80767084",
    69 => x"05580871",
    70 => x"5e5e577c",
    71 => x"7084055e",
    72 => x"0858805b",
    73 => x"77982a78",
    74 => x"882b5953",
    75 => x"72893876",
    76 => x"5e848080",
    77 => x"84bc047b",
    78 => x"802e81d8",
    79 => x"38805c72",
    80 => x"80e42ea1",
    81 => x"387280e4",
    82 => x"268e3872",
    83 => x"80e32e80",
    84 => x"f5388480",
    85 => x"8083d404",
    86 => x"7280f32e",
    87 => x"80d03884",
    88 => x"808083d4",
    89 => x"04758417",
    90 => x"71087e5c",
    91 => x"56575287",
    92 => x"55739c2a",
    93 => x"74842b55",
    94 => x"5271802e",
    95 => x"83388159",
    96 => x"8972258a",
    97 => x"38b71252",
    98 => x"84808083",
    99 => x"9104b012",
   100 => x"5278802e",
   101 => x"89387151",
   102 => x"84808081",
   103 => x"842dff15",
   104 => x"55748025",
   105 => x"cc388054",
   106 => x"84808083",
   107 => x"ed047584",
   108 => x"17710870",
   109 => x"545c5752",
   110 => x"84808081",
   111 => x"ab2d7b54",
   112 => x"84808083",
   113 => x"ed047584",
   114 => x"17710855",
   115 => x"57528480",
   116 => x"8084a404",
   117 => x"a5518480",
   118 => x"8081842d",
   119 => x"72518480",
   120 => x"8081842d",
   121 => x"82175784",
   122 => x"808084af",
   123 => x"0473ff15",
   124 => x"55528072",
   125 => x"25b93879",
   126 => x"7081055b",
   127 => x"84808080",
   128 => x"af2d7052",
   129 => x"53848080",
   130 => x"81842d81",
   131 => x"17578480",
   132 => x"8083ed04",
   133 => x"72a52e09",
   134 => x"81068938",
   135 => x"815c8480",
   136 => x"8084af04",
   137 => x"72518480",
   138 => x"8081842d",
   139 => x"81175781",
   140 => x"1b5b837b",
   141 => x"25fded38",
   142 => x"72fde038",
   143 => x"7d848080",
   144 => x"93900c02",
   145 => x"bc050d04",
   146 => x"02f4050d",
   147 => x"74765253",
   148 => x"80712590",
   149 => x"38705272",
   150 => x"70840554",
   151 => x"08ff1353",
   152 => x"5171f438",
   153 => x"028c050d",
   154 => x"0402d805",
   155 => x"0d7b7d5b",
   156 => x"56810b84",
   157 => x"80808d94",
   158 => x"59578359",
   159 => x"7708760c",
   160 => x"75087808",
   161 => x"56547375",
   162 => x"2e943875",
   163 => x"08537452",
   164 => x"8480808d",
   165 => x"a4518480",
   166 => x"8082812d",
   167 => x"80577952",
   168 => x"75518480",
   169 => x"8084c82d",
   170 => x"75085473",
   171 => x"752e9438",
   172 => x"75085374",
   173 => x"52848080",
   174 => x"8de45184",
   175 => x"80808281",
   176 => x"2d8057ff",
   177 => x"19841959",
   178 => x"59788025",
   179 => x"ffae3876",
   180 => x"84808093",
   181 => x"900c02a8",
   182 => x"050d0402",
   183 => x"ec050d76",
   184 => x"54815585",
   185 => x"aad5aad5",
   186 => x"740cfad5",
   187 => x"aad5aa0b",
   188 => x"8c150ccc",
   189 => x"74848080",
   190 => x"80c42db3",
   191 => x"0b8f1584",
   192 => x"808080c4",
   193 => x"2d730853",
   194 => x"72fce2d5",
   195 => x"aad52e92",
   196 => x"38730852",
   197 => x"8480808e",
   198 => x"a4518480",
   199 => x"8082812d",
   200 => x"80558c14",
   201 => x"085372fa",
   202 => x"d5aad4b3",
   203 => x"2e93388c",
   204 => x"14085284",
   205 => x"80808ee0",
   206 => x"51848080",
   207 => x"82812d80",
   208 => x"55775273",
   209 => x"51848080",
   210 => x"84c82d73",
   211 => x"085372fc",
   212 => x"e2d5aad5",
   213 => x"2e923873",
   214 => x"08528480",
   215 => x"808f9c51",
   216 => x"84808082",
   217 => x"812d8055",
   218 => x"8c140853",
   219 => x"72fad5aa",
   220 => x"d4b32e93",
   221 => x"388c1408",
   222 => x"52848080",
   223 => x"8fd85184",
   224 => x"80808281",
   225 => x"2d805574",
   226 => x"84808093",
   227 => x"900c0294",
   228 => x"050d0402",
   229 => x"c4050d60",
   230 => x"5e806290",
   231 => x"808029ff",
   232 => x"05848080",
   233 => x"9094535e",
   234 => x"5c848080",
   235 => x"82812d80",
   236 => x"e1b35780",
   237 => x"fe5bae51",
   238 => x"84808081",
   239 => x"842d7610",
   240 => x"70962a70",
   241 => x"81065156",
   242 => x"5774802e",
   243 => x"85387681",
   244 => x"07577695",
   245 => x"2a708106",
   246 => x"51557480",
   247 => x"2e853876",
   248 => x"81325778",
   249 => x"77077d06",
   250 => x"775b598f",
   251 => x"ffff5876",
   252 => x"bfffff06",
   253 => x"707a3282",
   254 => x"2b7f1151",
   255 => x"57760c76",
   256 => x"1070962a",
   257 => x"70810651",
   258 => x"56577480",
   259 => x"2e853876",
   260 => x"81075776",
   261 => x"952a7081",
   262 => x"06515574",
   263 => x"802e8538",
   264 => x"76813257",
   265 => x"ff185877",
   266 => x"8025c438",
   267 => x"79578fff",
   268 => x"ff5876bf",
   269 => x"ffff0670",
   270 => x"7a32822b",
   271 => x"7f117008",
   272 => x"51515656",
   273 => x"74762eab",
   274 => x"38807c53",
   275 => x"84808090",
   276 => x"a4525f84",
   277 => x"80808281",
   278 => x"2d745475",
   279 => x"53755284",
   280 => x"808090b8",
   281 => x"51848080",
   282 => x"82812d7e",
   283 => x"5c848080",
   284 => x"88f60481",
   285 => x"1c5c7610",
   286 => x"70962a70",
   287 => x"81065156",
   288 => x"5774802e",
   289 => x"85387681",
   290 => x"07577695",
   291 => x"2a708106",
   292 => x"51557480",
   293 => x"2e853876",
   294 => x"813257ff",
   295 => x"18587780",
   296 => x"25ff8f38",
   297 => x"ff1b5b7a",
   298 => x"fe8c388a",
   299 => x"51848080",
   300 => x"81842d7e",
   301 => x"84808093",
   302 => x"900c02bc",
   303 => x"050d0402",
   304 => x"d0050d7d",
   305 => x"5b815a80",
   306 => x"5980c07a",
   307 => x"595c85ad",
   308 => x"a989bb7b",
   309 => x"0c795781",
   310 => x"56975577",
   311 => x"7607822b",
   312 => x"7b115154",
   313 => x"85ada989",
   314 => x"bb740c75",
   315 => x"10ff1656",
   316 => x"56748025",
   317 => x"e6387710",
   318 => x"81185858",
   319 => x"987725d7",
   320 => x"387e527a",
   321 => x"51848080",
   322 => x"84c82d81",
   323 => x"58ff8787",
   324 => x"a5c37b0c",
   325 => x"97577782",
   326 => x"2b7b1170",
   327 => x"08565656",
   328 => x"73ff8787",
   329 => x"a5c32e09",
   330 => x"81068b38",
   331 => x"78780759",
   332 => x"8480808a",
   333 => x"d5047408",
   334 => x"547385ad",
   335 => x"a989bb2e",
   336 => x"94388075",
   337 => x"08547653",
   338 => x"84808090",
   339 => x"e0525a84",
   340 => x"80808281",
   341 => x"2d7710ff",
   342 => x"18585876",
   343 => x"8025ffb6",
   344 => x"3878822b",
   345 => x"5978802e",
   346 => x"80e33878",
   347 => x"52848080",
   348 => x"91805184",
   349 => x"80808281",
   350 => x"2d78992a",
   351 => x"81327081",
   352 => x"06700981",
   353 => x"05707207",
   354 => x"7009709f",
   355 => x"2c7f067e",
   356 => x"109fffff",
   357 => x"fe066281",
   358 => x"2a435f5f",
   359 => x"51515651",
   360 => x"5578d638",
   361 => x"79098105",
   362 => x"707b079f",
   363 => x"2a51547b",
   364 => x"bf269838",
   365 => x"73802e93",
   366 => x"38848080",
   367 => x"91985184",
   368 => x"80808281",
   369 => x"2d848080",
   370 => x"8bcd0481",
   371 => x"5c7b5284",
   372 => x"808091e4",
   373 => x"51848080",
   374 => x"82812d7b",
   375 => x"84808093",
   376 => x"900c02b0",
   377 => x"050d0402",
   378 => x"f4050d88",
   379 => x"bd0bff88",
   380 => x"0ca08052",
   381 => x"80518480",
   382 => x"8084e92d",
   383 => x"84808093",
   384 => x"9008802e",
   385 => x"8d388480",
   386 => x"8092a051",
   387 => x"84808082",
   388 => x"812da080",
   389 => x"52805184",
   390 => x"808085db",
   391 => x"2d848080",
   392 => x"93900880",
   393 => x"2e8d3884",
   394 => x"808092c4",
   395 => x"51848080",
   396 => x"82812da0",
   397 => x"80528051",
   398 => x"84808089",
   399 => x"bf2d8480",
   400 => x"80939008",
   401 => x"53848080",
   402 => x"93900880",
   403 => x"2e8d3884",
   404 => x"808092e0",
   405 => x"51848080",
   406 => x"82812d72",
   407 => x"52805184",
   408 => x"80808793",
   409 => x"2d848080",
   410 => x"93900880",
   411 => x"2eff8238",
   412 => x"84808092",
   413 => x"f8518480",
   414 => x"8082812d",
   415 => x"8480808b",
   416 => x"f1040000",
   417 => x"00ffffff",
   418 => x"ff00ffff",
   419 => x"ffff00ff",
   420 => x"ffffff00",
   421 => x"00000000",
   422 => x"55555555",
   423 => x"aaaaaaaa",
   424 => x"ffffffff",
   425 => x"53616e69",
   426 => x"74792063",
   427 => x"6865636b",
   428 => x"20666169",
   429 => x"6c656420",
   430 => x"28626566",
   431 => x"6f726520",
   432 => x"63616368",
   433 => x"65207265",
   434 => x"66726573",
   435 => x"6829206f",
   436 => x"6e203078",
   437 => x"25642028",
   438 => x"676f7420",
   439 => x"30782564",
   440 => x"290a0000",
   441 => x"53616e69",
   442 => x"74792063",
   443 => x"6865636b",
   444 => x"20666169",
   445 => x"6c656420",
   446 => x"28616674",
   447 => x"65722063",
   448 => x"61636865",
   449 => x"20726566",
   450 => x"72657368",
   451 => x"29206f6e",
   452 => x"20307825",
   453 => x"64202867",
   454 => x"6f742030",
   455 => x"78256429",
   456 => x"0a000000",
   457 => x"42797465",
   458 => x"20636865",
   459 => x"636b2066",
   460 => x"61696c65",
   461 => x"64202862",
   462 => x"65666f72",
   463 => x"65206361",
   464 => x"63686520",
   465 => x"72656672",
   466 => x"65736829",
   467 => x"20617420",
   468 => x"30202867",
   469 => x"6f742030",
   470 => x"78256429",
   471 => x"0a000000",
   472 => x"42797465",
   473 => x"20636865",
   474 => x"636b2066",
   475 => x"61696c65",
   476 => x"64202862",
   477 => x"65666f72",
   478 => x"65206361",
   479 => x"63686520",
   480 => x"72656672",
   481 => x"65736829",
   482 => x"20617420",
   483 => x"33202867",
   484 => x"6f742030",
   485 => x"78256429",
   486 => x"0a000000",
   487 => x"42797465",
   488 => x"20636865",
   489 => x"636b2066",
   490 => x"61696c65",
   491 => x"64202861",
   492 => x"66746572",
   493 => x"20636163",
   494 => x"68652072",
   495 => x"65667265",
   496 => x"73682920",
   497 => x"61742030",
   498 => x"2028676f",
   499 => x"74203078",
   500 => x"2564290a",
   501 => x"00000000",
   502 => x"42797465",
   503 => x"20636865",
   504 => x"636b2066",
   505 => x"61696c65",
   506 => x"64202861",
   507 => x"66746572",
   508 => x"20636163",
   509 => x"68652072",
   510 => x"65667265",
   511 => x"73682920",
   512 => x"61742033",
   513 => x"2028676f",
   514 => x"74203078",
   515 => x"2564290a",
   516 => x"00000000",
   517 => x"43686563",
   518 => x"6b696e67",
   519 => x"206d656d",
   520 => x"6f727900",
   521 => x"30782564",
   522 => x"20676f6f",
   523 => x"64207265",
   524 => x"6164732c",
   525 => x"20000000",
   526 => x"4572726f",
   527 => x"72206174",
   528 => x"20307825",
   529 => x"642c2065",
   530 => x"78706563",
   531 => x"74656420",
   532 => x"30782564",
   533 => x"2c20676f",
   534 => x"74203078",
   535 => x"25640a00",
   536 => x"42616420",
   537 => x"64617461",
   538 => x"20666f75",
   539 => x"6e642061",
   540 => x"74203078",
   541 => x"25642028",
   542 => x"30782564",
   543 => x"290a0000",
   544 => x"416c6961",
   545 => x"73657320",
   546 => x"666f756e",
   547 => x"64206174",
   548 => x"20307825",
   549 => x"640a0000",
   550 => x"28416c69",
   551 => x"61736573",
   552 => x"2070726f",
   553 => x"6261626c",
   554 => x"79207369",
   555 => x"6d706c79",
   556 => x"20696e64",
   557 => x"69636174",
   558 => x"65207468",
   559 => x"61742052",
   560 => x"414d0a69",
   561 => x"7320736d",
   562 => x"616c6c65",
   563 => x"72207468",
   564 => x"616e2036",
   565 => x"34206d65",
   566 => x"67616279",
   567 => x"74657329",
   568 => x"0a000000",
   569 => x"53445241",
   570 => x"4d207369",
   571 => x"7a652028",
   572 => x"61737375",
   573 => x"6d696e67",
   574 => x"206e6f20",
   575 => x"61646472",
   576 => x"65737320",
   577 => x"6661756c",
   578 => x"74732920",
   579 => x"69732030",
   580 => x"78256420",
   581 => x"6d656761",
   582 => x"62797465",
   583 => x"730a0000",
   584 => x"46697273",
   585 => x"74207374",
   586 => x"61676520",
   587 => x"73616e69",
   588 => x"74792063",
   589 => x"6865636b",
   590 => x"20706173",
   591 => x"7365642e",
   592 => x"0a000000",
   593 => x"42797465",
   594 => x"20286471",
   595 => x"6d292063",
   596 => x"6865636b",
   597 => x"20706173",
   598 => x"7365640a",
   599 => x"00000000",
   600 => x"41646472",
   601 => x"65737320",
   602 => x"63686563",
   603 => x"6b207061",
   604 => x"73736564",
   605 => x"2e0a0000",
   606 => x"4c465352",
   607 => x"20636865",
   608 => x"636b2070",
   609 => x"61737365",
   610 => x"642e0a0a",
   611 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

