-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity SDRAMTest_ROM is
generic
	(
		maxAddrBit : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end SDRAMTest_ROM;

architecture arch of SDRAMTest_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBit+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0ba08080",
     1 => x"df040000",
     2 => x"80047004",
     3 => x"71fd0608",
     4 => x"72830609",
     5 => x"81058205",
     6 => x"832b2a83",
     7 => x"ffff0652",
     8 => x"0471fc06",
     9 => x"08728306",
    10 => x"09810583",
    11 => x"05101010",
    12 => x"2a81ff06",
    13 => x"520471fc",
    14 => x"06080ba0",
    15 => x"808ca073",
    16 => x"83061010",
    17 => x"05080673",
    18 => x"81ff0673",
    19 => x"83060981",
    20 => x"05830510",
    21 => x"10102b07",
    22 => x"72fc060c",
    23 => x"5151040b",
    24 => x"a08080ea",
    25 => x"0ba0808b",
    26 => x"96040ba0",
    27 => x"8080ea04",
    28 => x"00000002",
    29 => x"f8050d73",
    30 => x"52ff8408",
    31 => x"70882a70",
    32 => x"81065151",
    33 => x"5170802e",
    34 => x"f03871ff",
    35 => x"840c71a0",
    36 => x"8092ac0c",
    37 => x"0288050d",
    38 => x"0402f005",
    39 => x"0d755380",
    40 => x"73a08080",
    41 => x"a12d7081",
    42 => x"ff065353",
    43 => x"5470742e",
    44 => x"b0387181",
    45 => x"ff068114",
    46 => x"5452ff84",
    47 => x"0870882a",
    48 => x"70810651",
    49 => x"51517080",
    50 => x"2ef03871",
    51 => x"ff840c81",
    52 => x"1473a080",
    53 => x"80a12d70",
    54 => x"81ff0653",
    55 => x"535470d2",
    56 => x"3873a080",
    57 => x"92ac0c02",
    58 => x"90050d04",
    59 => x"02c4050d",
    60 => x"0280c005",
    61 => x"a080938c",
    62 => x"5b568076",
    63 => x"70840558",
    64 => x"08715e5e",
    65 => x"577c7084",
    66 => x"055e0858",
    67 => x"805b7798",
    68 => x"2a78882b",
    69 => x"59537288",
    70 => x"38765ea0",
    71 => x"80849504",
    72 => x"7b802e81",
    73 => x"ca38805c",
    74 => x"7280e42e",
    75 => x"9f387280",
    76 => x"e4268d38",
    77 => x"7280e32e",
    78 => x"80ee38a0",
    79 => x"8083b504",
    80 => x"7280f32e",
    81 => x"80cc38a0",
    82 => x"8083b504",
    83 => x"75841771",
    84 => x"087e5c56",
    85 => x"57528755",
    86 => x"739c2a74",
    87 => x"842b5552",
    88 => x"71802e83",
    89 => x"38815989",
    90 => x"72258938",
    91 => x"b71252a0",
    92 => x"8082f704",
    93 => x"b0125278",
    94 => x"802e8838",
    95 => x"7151a080",
    96 => x"80f32dff",
    97 => x"15557480",
    98 => x"25ce3880",
    99 => x"54a08083",
   100 => x"cb047584",
   101 => x"17710870",
   102 => x"545c5752",
   103 => x"a0808199",
   104 => x"2d7b54a0",
   105 => x"8083cb04",
   106 => x"75841771",
   107 => x"08555752",
   108 => x"a08083fe",
   109 => x"04a551a0",
   110 => x"8080f32d",
   111 => x"7251a080",
   112 => x"80f32d82",
   113 => x"1757a080",
   114 => x"84880473",
   115 => x"ff155552",
   116 => x"807225b4",
   117 => x"38797081",
   118 => x"055ba080",
   119 => x"80a12d70",
   120 => x"5253a080",
   121 => x"80f32d81",
   122 => x"1757a080",
   123 => x"83cb0472",
   124 => x"a52e0981",
   125 => x"06883881",
   126 => x"5ca08084",
   127 => x"88047251",
   128 => x"a08080f3",
   129 => x"2d811757",
   130 => x"811b5b83",
   131 => x"7b25fdfe",
   132 => x"3872fdf1",
   133 => x"387da080",
   134 => x"92ac0c02",
   135 => x"bc050d04",
   136 => x"02f4050d",
   137 => x"74765253",
   138 => x"80712590",
   139 => x"38705272",
   140 => x"70840554",
   141 => x"08ff1353",
   142 => x"5171f438",
   143 => x"028c050d",
   144 => x"0402d805",
   145 => x"0d7b7d5b",
   146 => x"56810ba0",
   147 => x"808cb059",
   148 => x"57835977",
   149 => x"08760c75",
   150 => x"08780856",
   151 => x"5473752e",
   152 => x"92387508",
   153 => x"537452a0",
   154 => x"808cc051",
   155 => x"a08081ec",
   156 => x"2d805779",
   157 => x"527551a0",
   158 => x"8084a02d",
   159 => x"75085473",
   160 => x"752e9238",
   161 => x"75085374",
   162 => x"52a0808d",
   163 => x"8051a080",
   164 => x"81ec2d80",
   165 => x"57ff1984",
   166 => x"19595978",
   167 => x"8025ffb3",
   168 => x"3876a080",
   169 => x"92ac0c02",
   170 => x"a8050d04",
   171 => x"02ec050d",
   172 => x"76548155",
   173 => x"85aad5aa",
   174 => x"d5740cfa",
   175 => x"d5aad5aa",
   176 => x"0b8c150c",
   177 => x"cc74a080",
   178 => x"80b62db3",
   179 => x"0b8f15a0",
   180 => x"8080b62d",
   181 => x"73085372",
   182 => x"fce2d5aa",
   183 => x"d52e9038",
   184 => x"730852a0",
   185 => x"808dc051",
   186 => x"a08081ec",
   187 => x"2d80558c",
   188 => x"14085372",
   189 => x"fad5aad4",
   190 => x"b32e9138",
   191 => x"8c140852",
   192 => x"a0808dfc",
   193 => x"51a08081",
   194 => x"ec2d8055",
   195 => x"77527351",
   196 => x"a08084a0",
   197 => x"2d730853",
   198 => x"72fce2d5",
   199 => x"aad52e90",
   200 => x"38730852",
   201 => x"a0808eb8",
   202 => x"51a08081",
   203 => x"ec2d8055",
   204 => x"8c140853",
   205 => x"72fad5aa",
   206 => x"d4b32e91",
   207 => x"388c1408",
   208 => x"52a0808e",
   209 => x"f451a080",
   210 => x"81ec2d80",
   211 => x"5574a080",
   212 => x"92ac0c02",
   213 => x"94050d04",
   214 => x"02c4050d",
   215 => x"605e8062",
   216 => x"90808029",
   217 => x"ff05a080",
   218 => x"8fb0535e",
   219 => x"5ca08081",
   220 => x"ec2d80e1",
   221 => x"b35780fe",
   222 => x"5bae51a0",
   223 => x"8080f32d",
   224 => x"76107096",
   225 => x"2a708106",
   226 => x"51565774",
   227 => x"802e8538",
   228 => x"76810757",
   229 => x"76952a70",
   230 => x"81065155",
   231 => x"74802e85",
   232 => x"38768132",
   233 => x"57787707",
   234 => x"7d06775b",
   235 => x"598fffff",
   236 => x"5876bfff",
   237 => x"ff06707a",
   238 => x"32822b7f",
   239 => x"11515776",
   240 => x"0c761070",
   241 => x"962a7081",
   242 => x"06515657",
   243 => x"74802e85",
   244 => x"38768107",
   245 => x"5776952a",
   246 => x"70810651",
   247 => x"5574802e",
   248 => x"85387681",
   249 => x"3257ff18",
   250 => x"58778025",
   251 => x"c4387957",
   252 => x"8fffff58",
   253 => x"76bfffff",
   254 => x"06707a32",
   255 => x"822b7f11",
   256 => x"70085151",
   257 => x"56567476",
   258 => x"2ea63880",
   259 => x"7c53a080",
   260 => x"8fc0525f",
   261 => x"a08081ec",
   262 => x"2d745475",
   263 => x"537552a0",
   264 => x"808fd451",
   265 => x"a08081ec",
   266 => x"2d7e5ca0",
   267 => x"8088b304",
   268 => x"811c5c76",
   269 => x"1070962a",
   270 => x"70810651",
   271 => x"56577480",
   272 => x"2e853876",
   273 => x"81075776",
   274 => x"952a7081",
   275 => x"06515574",
   276 => x"802e8538",
   277 => x"76813257",
   278 => x"ff185877",
   279 => x"8025ff94",
   280 => x"38ff1b5b",
   281 => x"7afe9238",
   282 => x"8a51a080",
   283 => x"80f32d7e",
   284 => x"a08092ac",
   285 => x"0c02bc05",
   286 => x"0d0402d0",
   287 => x"050d7d5b",
   288 => x"815a8059",
   289 => x"80c07a59",
   290 => x"5c85ada9",
   291 => x"89bb7b0c",
   292 => x"79578156",
   293 => x"97557776",
   294 => x"07822b7b",
   295 => x"11515485",
   296 => x"ada989bb",
   297 => x"740c7510",
   298 => x"ff165656",
   299 => x"748025e6",
   300 => x"38771081",
   301 => x"18585898",
   302 => x"7725d738",
   303 => x"7e527a51",
   304 => x"a08084a0",
   305 => x"2d8158ff",
   306 => x"8787a5c3",
   307 => x"7b0c9757",
   308 => x"77822b7b",
   309 => x"11700856",
   310 => x"565673ff",
   311 => x"8787a5c3",
   312 => x"2e098106",
   313 => x"8a387878",
   314 => x"0759a080",
   315 => x"8a8c0474",
   316 => x"08547385",
   317 => x"ada989bb",
   318 => x"2e923880",
   319 => x"75085476",
   320 => x"53a0808f",
   321 => x"fc525aa0",
   322 => x"8081ec2d",
   323 => x"7710ff18",
   324 => x"58587680",
   325 => x"25ffb938",
   326 => x"78822b59",
   327 => x"78802e80",
   328 => x"de387852",
   329 => x"a080909c",
   330 => x"51a08081",
   331 => x"ec2d7899",
   332 => x"2a813270",
   333 => x"81067009",
   334 => x"81057072",
   335 => x"07700970",
   336 => x"9f2c7f06",
   337 => x"7e109fff",
   338 => x"fffe0662",
   339 => x"812a435f",
   340 => x"5f515156",
   341 => x"515578d6",
   342 => x"38790981",
   343 => x"05707b07",
   344 => x"9f2a5154",
   345 => x"7bbf2695",
   346 => x"3873802e",
   347 => x"9038a080",
   348 => x"90b451a0",
   349 => x"8081ec2d",
   350 => x"a0808aff",
   351 => x"04815c7b",
   352 => x"52a08091",
   353 => x"8051a080",
   354 => x"81ec2d7b",
   355 => x"a08092ac",
   356 => x"0c02b005",
   357 => x"0d0402f4",
   358 => x"050d88bd",
   359 => x"0bff880c",
   360 => x"a0805280",
   361 => x"51a08084",
   362 => x"c12da080",
   363 => x"92ac0880",
   364 => x"2e8b38a0",
   365 => x"8091bc51",
   366 => x"a08081ec",
   367 => x"2da08052",
   368 => x"8051a080",
   369 => x"85ac2da0",
   370 => x"8092ac08",
   371 => x"802e8b38",
   372 => x"a08091e0",
   373 => x"51a08081",
   374 => x"ec2da080",
   375 => x"528051a0",
   376 => x"8088fa2d",
   377 => x"a08092ac",
   378 => x"0853a080",
   379 => x"92ac0880",
   380 => x"2e8b38a0",
   381 => x"8091fc51",
   382 => x"a08081ec",
   383 => x"2d725280",
   384 => x"51a08086",
   385 => x"d82da080",
   386 => x"92ac0880",
   387 => x"2eff9138",
   388 => x"a0809294",
   389 => x"51a08081",
   390 => x"ec2da080",
   391 => x"8ba00400",
   392 => x"00ffffff",
   393 => x"ff00ffff",
   394 => x"ffff00ff",
   395 => x"ffffff00",
   396 => x"00000000",
   397 => x"55555555",
   398 => x"aaaaaaaa",
   399 => x"ffffffff",
   400 => x"53616e69",
   401 => x"74792063",
   402 => x"6865636b",
   403 => x"20666169",
   404 => x"6c656420",
   405 => x"28626566",
   406 => x"6f726520",
   407 => x"63616368",
   408 => x"65207265",
   409 => x"66726573",
   410 => x"6829206f",
   411 => x"6e203078",
   412 => x"25642028",
   413 => x"676f7420",
   414 => x"30782564",
   415 => x"290a0000",
   416 => x"53616e69",
   417 => x"74792063",
   418 => x"6865636b",
   419 => x"20666169",
   420 => x"6c656420",
   421 => x"28616674",
   422 => x"65722063",
   423 => x"61636865",
   424 => x"20726566",
   425 => x"72657368",
   426 => x"29206f6e",
   427 => x"20307825",
   428 => x"64202867",
   429 => x"6f742030",
   430 => x"78256429",
   431 => x"0a000000",
   432 => x"42797465",
   433 => x"20636865",
   434 => x"636b2066",
   435 => x"61696c65",
   436 => x"64202862",
   437 => x"65666f72",
   438 => x"65206361",
   439 => x"63686520",
   440 => x"72656672",
   441 => x"65736829",
   442 => x"20617420",
   443 => x"30202867",
   444 => x"6f742030",
   445 => x"78256429",
   446 => x"0a000000",
   447 => x"42797465",
   448 => x"20636865",
   449 => x"636b2066",
   450 => x"61696c65",
   451 => x"64202862",
   452 => x"65666f72",
   453 => x"65206361",
   454 => x"63686520",
   455 => x"72656672",
   456 => x"65736829",
   457 => x"20617420",
   458 => x"33202867",
   459 => x"6f742030",
   460 => x"78256429",
   461 => x"0a000000",
   462 => x"42797465",
   463 => x"20636865",
   464 => x"636b2066",
   465 => x"61696c65",
   466 => x"64202861",
   467 => x"66746572",
   468 => x"20636163",
   469 => x"68652072",
   470 => x"65667265",
   471 => x"73682920",
   472 => x"61742030",
   473 => x"2028676f",
   474 => x"74203078",
   475 => x"2564290a",
   476 => x"00000000",
   477 => x"42797465",
   478 => x"20636865",
   479 => x"636b2066",
   480 => x"61696c65",
   481 => x"64202861",
   482 => x"66746572",
   483 => x"20636163",
   484 => x"68652072",
   485 => x"65667265",
   486 => x"73682920",
   487 => x"61742033",
   488 => x"2028676f",
   489 => x"74203078",
   490 => x"2564290a",
   491 => x"00000000",
   492 => x"43686563",
   493 => x"6b696e67",
   494 => x"206d656d",
   495 => x"6f727900",
   496 => x"30782564",
   497 => x"20676f6f",
   498 => x"64207265",
   499 => x"6164732c",
   500 => x"20000000",
   501 => x"4572726f",
   502 => x"72206174",
   503 => x"20307825",
   504 => x"642c2065",
   505 => x"78706563",
   506 => x"74656420",
   507 => x"30782564",
   508 => x"2c20676f",
   509 => x"74203078",
   510 => x"25640a00",
   511 => x"42616420",
   512 => x"64617461",
   513 => x"20666f75",
   514 => x"6e642061",
   515 => x"74203078",
   516 => x"25642028",
   517 => x"30782564",
   518 => x"290a0000",
   519 => x"416c6961",
   520 => x"73657320",
   521 => x"666f756e",
   522 => x"64206174",
   523 => x"20307825",
   524 => x"640a0000",
   525 => x"28416c69",
   526 => x"61736573",
   527 => x"2070726f",
   528 => x"6261626c",
   529 => x"79207369",
   530 => x"6d706c79",
   531 => x"20696e64",
   532 => x"69636174",
   533 => x"65207468",
   534 => x"61742052",
   535 => x"414d0a69",
   536 => x"7320736d",
   537 => x"616c6c65",
   538 => x"72207468",
   539 => x"616e2036",
   540 => x"34206d65",
   541 => x"67616279",
   542 => x"74657329",
   543 => x"0a000000",
   544 => x"53445241",
   545 => x"4d207369",
   546 => x"7a652028",
   547 => x"61737375",
   548 => x"6d696e67",
   549 => x"206e6f20",
   550 => x"61646472",
   551 => x"65737320",
   552 => x"6661756c",
   553 => x"74732920",
   554 => x"69732030",
   555 => x"78256420",
   556 => x"6d656761",
   557 => x"62797465",
   558 => x"730a0000",
   559 => x"46697273",
   560 => x"74207374",
   561 => x"61676520",
   562 => x"73616e69",
   563 => x"74792063",
   564 => x"6865636b",
   565 => x"20706173",
   566 => x"7365642e",
   567 => x"0a000000",
   568 => x"42797465",
   569 => x"20286471",
   570 => x"6d292063",
   571 => x"6865636b",
   572 => x"20706173",
   573 => x"7365640a",
   574 => x"00000000",
   575 => x"41646472",
   576 => x"65737320",
   577 => x"63686563",
   578 => x"6b207061",
   579 => x"73736564",
   580 => x"2e0a0000",
   581 => x"4c465352",
   582 => x"20636865",
   583 => x"636b2070",
   584 => x"61737365",
   585 => x"642e0a0a",
   586 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBit downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBit downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBit downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBit downto 2))));
		end if;
	end if;
end process;


end arch;

